library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity waveform_generator is 

end;

architecture behavioural of waveform_generator is

begin

end;
