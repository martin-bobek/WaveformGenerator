library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tb_waveform_generator is end;

architecture Behavioral of tb_waveform_generator is
    component waveform_generator is 
    end component;
begin


end Behavioral;
